interface intf(input logic clk,reset);
  logic valid;
  logic a,b;
  logic sum,carry;
endinterface